../microcontroller/microcontroller.vhd