../Alu/memory_cell.vhd