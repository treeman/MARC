../Alu/Memory_Cell_DualPort.vhd