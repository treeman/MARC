../Alu/ALU.vhd